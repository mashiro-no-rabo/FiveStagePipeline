`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:        Team.TeaWhen
// Engineer:       AquarHEAD L.
// 
// Create Date:    21:27:58 04/25/2013 
// Design Name: 
// Header Name:    ALUOP 
// Project Name:   Five Stage Pipeline CPU
// Target Devices: Spartan3E Starter Kit
// Tool versions:  Xilinx ISE 14.1
// Description:    I love @Lilian_Ye
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

//ALU CODE
`define ALU_ADD 4'b0000
`define ALU_SUB 4'b0010
`define ALU_AND 4'b0100
`define ALU_OR  4'b0101
`define ALU_NOR 4'b0111
`define ALU_SLT 4'b1000
`define ALU_SLL 4'b1100
`define ALU_SRL 4'b1101
`define ALU_SRA 4'b1111
//`define ALU_NONE 4'b1110
